library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity; cat
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity; cat
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity; cat
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity; cat
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity; cat
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity; cat
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity;
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity;
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity;
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity;
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity;
library ieee;
use ieee.std_logic_1164.all;

entity test_tb is



end entity;
